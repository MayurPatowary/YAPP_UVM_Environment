module hw_top;

  // Clock and reset signals
  logic [31:0]  clock_period;
  logic         run_clock;
  logic         clock;
  logic         reset;

  // YAPP Interface to the DUT
  yapp_if in0(clock, reset);

  // Clock and Reset Interface to the DUT
  clock_and_reset_if cr0(clock, reset, run_clock, clock_period);
  // clock_and_reset_if interface doesn't generate clk signal directly but supplies control signals (run_clock and clock_period) to the clkgen instance. The clkgen 
  // generates the clk and the clk is passed back into clock_and_reset_if to synchronize the reset generation. 
  // These control signals are generated by the interface when sequences execute on Clock and Reset UVC.
  // So, the clock and reset interface has a clock input port but reset, run clock, and clock period output ports.

  // HBUS Interface to the DUT
  hbus_if hb0(clock, reset);

   // Channel Interfaces to the DUT
   channel_if ch0(clock, reset);
   channel_if ch1(clock, reset);
   channel_if ch2(clock, reset);

  // CLKGEN module generates clock
  clkgen clkgen (
    .clock(clock),
    .run_clock(run_clock),
    .clock_period(clock_period)
  );
  // The run clock and clock period interface outputs are connected to the clkgen ports. This allows Clock and Reset UVC sequences to control the clock generation.

  yapp_router dut(
    .reset(reset),
    .clock(clock),
    .error(),

    // YAPP interface
    .in_data(in0.in_data),
    .in_data_vld(in0.in_data_vld),
    .in_suspend(in0.in_suspend),

    // Output Channels
    //Channel 0
    .data_0(ch0.data),
    .data_vld_0(ch0.data_vld),
    .suspend_0(ch0.suspend),
    
    //Channel 1
    .data_1(ch1.data),
    .data_vld_1(ch1.data_vld),
    .suspend_1(ch1.suspend),
    
    //Channel 2
    .data_2(ch2.data),
    .data_vld_2(ch2.data_vld),
    .suspend_2(ch2.suspend),

    // HBUS Interface 
    .haddr(hb0.haddr),
    .hdata(hb0.hdata_w),
    .hen(hb0.hen),
    .hwr_rd(hb0.hwr_rd)
    );

endmodule
